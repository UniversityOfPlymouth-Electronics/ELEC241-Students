library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ELEC233_ALU is

	-- Type Declaration (optional)

	-- Subtype Declaration (optional)
	constant WORD_WIDTH : natural := 8;
	
	-- Constant Declaration (optional)

	-- Signal Declaration (optional)

	-- Component Declaration (optional)

end ELEC233_ALU;


package body ELEC233_ALU is

	-- Type Declaration (optional)

	-- Subtype Declaration (optional)

	-- Constant Declaration (optional)

	-- Function Declaration (optional)

	-- Function Body (optional)

	-- Procedure Declaration (optional)

	-- Procedure Body (optional)

end ELEC233_ALU;
